LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY EK_TB IS END ENTITY;

ARCHITECTURE ARCH_EK_TB OF EK_TB IS
	COMPONENT EK IS PORT
	(
		CLK :  IN  STD_LOGIC;
		INIT :  IN  STD_LOGIC;
		RUN :  IN  STD_LOGIC;
		KEY :  IN  STD_LOGIC_VECTOR(127 DOWNTO 0);
		STATE_IN :  IN  STD_LOGIC_VECTOR(127 DOWNTO 0);
		STATE_OUT :  OUT  STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
	END COMPONENT;

	SIGNAL CLK :    STD_LOGIC := '0';
	SIGNAL INIT :    STD_LOGIC := '0';
	SIGNAL RUN :    STD_LOGIC := '0';
	SIGNAL KEY :    STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	SIGNAL STATE_IN :    STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	SIGNAL STATE_OUT :   STD_LOGIC_VECTOR(127 DOWNTO 0) := (OTHERS => '0');
	
	SIGNAL CLKp :time := 40 ns;
BEGIN
	tb: EK PORT MAP (CLK, INIT, RUN, KEY, STATE_IN, STATE_OUT);

	PROCESS
	BEGIN
		CLK <= '0'; wait for CLKp / 2;
		CLK <= '1'; wait for CLKp / 2;
	END PROCESS;

	PROCESS
	BEGIN
		INIT <= '1'; RUN <= '0'; KEY <= X"00000000000000000000000000000000"; STATE_IN <= X"00000000000000000000000000000000"; wait for CLKp;
		INIT <= '0'; RUN <= '1'; KEY <= X"00112233445566778899AABBCCDDEEFF"; STATE_IN <= X"00000000000000000000000000000000"; wait for 50*CLKp;
		--INIT <= '0'; RUN <= '1'; KEY <= X"00000000000000000000000000000000"; STATE_IN <= X"00000000000000000000000000000000"; wait for CLKp;

		wait;
	END PROCESS;
END ARCHITECTURE;