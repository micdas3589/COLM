LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY KEY_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DATA_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		KEY		:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE ARCH_KEY_REG OF KEY_REG IS
	SIGNAL KEY_STATE	:STD_LOGIC_VECTOR(127 downto 0);
BEGIN
	PROCESS(CLK, INIT, KEY_STATE)
	BEGIN
		IF INIT = '1' THEN
			KEY_STATE	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				IF ADDR_WR = X"0" THEN
					KEY_STATE(127 downto 96)<= DATA_WR;
				END IF;
				IF ADDR_WR = X"1" THEN
					KEY_STATE(95 downto 64)	<= DATA_WR;
				END IF;
				IF ADDR_WR = X"2" THEN
					KEY_STATE(63 downto 32)	<= DATA_WR;
				END IF;
				IF ADDR_WR = X"3" THEN
					KEY_STATE(31 downto 0)	<= DATA_WR;
				END IF;
			END IF;
		END IF;
		
		KEY	<= KEY_STATE;
	END PROCESS;
END ARCHITECTURE;