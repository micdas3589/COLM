LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY ROUND_CTRL IS
	PORT (
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		RUN			:IN STD_LOGIC;
		LOAD_KEY		:OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE ROUND_CTRL_ARCH OF ROUND_CTRL IS
	SIGNAL LOADED_KEY	:STD_LOGIC := '0';
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			LOADED_KEY	<= '0';
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF RUN = '1' AND LOADED_KEY = '0' THEN
				LOADED_KEY	<= '1';
			END IF;
		END IF;
	END PROCESS;

	LOAD_KEY	<= '1'
					WHEN RUN = '1' AND LOADED_KEY = '0'
					ELSE '0';
END ARCHITECTURE;