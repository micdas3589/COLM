LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY CONTROL IS
	PORT (
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		WR				:IN STD_LOGIC;
		ADDR			:IN STD_LOGIC_VECTOR(31 downto 0);
		DRL_ASCD		:IN STD_LOGIC;
		DRL_PTX		:IN STD_LOGIC;
		WR_PTX		:OUT STD_LOGIC;
		WR_ASCD		:OUT STD_LOGIC;
		RD_PTX		:OUT STD_LOGIC;
		RD_ASCD		:OUT STD_LOGIC;
		RD_PARAMS	:OUT STD_LOGIC;
		WR_L			:OUT STD_LOGIC;
		DBL_L			:OUT STD_LOGIC;
		DBL_L1		:OUT STD_LOGIC;
		DBL_L2		:OUT STD_LOGIC;
		WR_IV			:OUT STD_LOGIC;
		RD_L			:OUT STD_LOGIC;
		RD_L1			:OUT STD_LOGIC;
		
		LOAD_KEY		:OUT STD_LOGIC;
		RUN_EK1		:OUT STD_LOGIC;
		RUN_EK2		:OUT STD_LOGIC;
		RUN_EK3		:OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE ARCH_CONTROL OF CONTROL IS
	SIGNAL COUNTER		:STD_LOGIC_VECTOR(15 downto 0);
	
	CONSTANT RUNNING	:STD_LOGIC := '1';
	CONSTANT IDLE		:STD_LOGIC := '0';
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			COUNTER	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF (WR = '1' AND ADDR = X"FFFFFFFF") OR COUNTER /= X"0" THEN
				IF COUNTER /= X"FFFF" THEN
					COUNTER	<= COUNTER + 1;
				END IF;
				IF COUNTER = X"0" THEN
					LOAD_KEY	<= '1'
				END IF;
				IF COUNTER <= X"2D" AND COUNTER <= X"59" AND DRL_ASCD = '1' THEN
					RUN_EK1	<= '1';
				END IF;
				IF COUNTER = X""
			END IF;
		END IF;
	END PROCESS;
	
	RUN_EK1		<= '1'
						WHEN COUNTER >= X"1" AND COUNTER <= X"2D"
						ELSE '0';
	WR_L			<= '1'
						WHEN COUNTER = X"2D" OR COUNTER = X"2E"
						ELSE '0';
	RD_PARAMS	<= '1'
						WHEN COUNTER = X"2F"
						ELSE '0';
	RD_L			<= '1'
						WHEN DRL_ASCD = '1'
						ELSE '0';
	RD_L1			<= '1'
						WHEN DRL_PTX = '1' AND DRL_ASCD = '0'
						ELSE '0';
	WR_PTX		<= '1'
						WHEN WR = '1' AND ADDR = X"11111111"
						ELSE '0';
	WR_ASCD		<= '1'
						WHEN WR = '1' AND ADDR = X"22222222"
						ELSE '0';
	LOAD_KEY		<= '1'
						WHEN COUNTER(1 downto 0) = X"1";
						ELSE '0';
END ARCHITECTURE;