LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY CONTROL IS
	PORT (
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		WR				:IN STD_LOGIC;
		RD				:IN STD_LOGIC;
		ADDR_WR		:IN STD_LOGIC_VECTOR(31 downto 0);
		DRL_ASCD		:IN STD_LOGIC;
		DRL_PTX		:IN STD_LOGIC;
		DRL_CTX		:IN STD_LOGIC;
		WR_PTX		:OUT STD_LOGIC;
		WR_ASCD		:OUT STD_LOGIC;
		WR_CTX		:OUT STD_LOGIC;
		RD_PTX		:OUT STD_LOGIC;
		RD_ASCD		:OUT STD_LOGIC;
		RD_PARAMS	:OUT STD_LOGIC;
		RD_CTX		:OUT STD_LOGIC;
		WR_L			:OUT STD_LOGIC;
		DBL_L			:OUT STD_LOGIC;
		DBL_L1		:OUT STD_LOGIC;
		DBL_L2		:OUT STD_LOGIC;
		WR_IV			:OUT STD_LOGIC;
		RD_L			:OUT STD_LOGIC;
		RD_L1			:OUT STD_LOGIC;
		WR_RO			:OUT STD_LOGIC;
		LOAD_IV		:OUT STD_LOGIC;
		INIT_EK1		:OUT STD_LOGIC;
		INIT_EK2		:OUT STD_LOGIC;
		INIT_EK3		:OUT STD_LOGIC;
		
		RUN_EK1		:OUT STD_LOGIC;
		RUN_EK2		:OUT STD_LOGIC;
		RUN_EK3		:OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE ARCH_CONTROL OF CONTROL IS
	SIGNAL COUNTER_ASCD	:STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL COUNTER_PTX	:STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL COUNTER_TAG	:STD_LOGIC_VECTOR(15 downto 0);
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			COUNTER_ASCD	<= (OTHERS => '0');
			COUNTER_PTX		<= (OTHERS => '0');
			COUNTER_TAG		<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF (WR = '1' AND ADDR_WR = X"FFFFFFFF") OR COUNTER_ASCD /= X"0" THEN
				IF COUNTER_ASCD /= X"8B" AND COUNTER_ASCD /= X"FF" THEN
					COUNTER_ASCD	<= COUNTER_ASCD + 1;
				END IF;
				IF COUNTER_ASCD = X"8B" THEN
					COUNTER_ASCD	<= X"5D";
				END IF;
				IF COUNTER_ASCD = X"8B" AND DRL_ASCD = '0' THEN
					COUNTER_ASCD	<= X"FF";
				END IF;
				
				IF COUNTER_ASCD = X"FF" AND COUNTER_PTX /= X"2F" AND COUNTER_PTX /= X"FF" THEN
					COUNTER_PTX	<= COUNTER_PTX + 1;
				END IF;
				IF COUNTER_PTX = X"2F" THEN
					COUNTER_PTX	<= X"01";
				END IF;
				IF COUNTER_PTX = X"2F" AND DRL_PTX = '0' THEN
					COUNTER_PTX	<= X"FF";
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	RUN_EK1		<= '1'
						WHEN (COUNTER_ASCD >= X"1" AND COUNTER_ASCD <= X"2E") -- GENERATE L
						  OR (COUNTER_ASCD >= X"30" AND COUNTER_ASCD <= X"5C") -- ENCRYPT PARAMS
						  OR (COUNTER_ASCD >= X"5E" AND COUNTER_ASCD <= X"8A") -- ENCRYPT ASCD
						  OR (COUNTER_PTX >= X"2" AND COUNTER_PTX <= X"2F") -- ENCRYPT PTX
						ELSE '0';
	INIT_EK1		<= '1'
						WHEN COUNTER_ASCD = X"00"
						  OR COUNTER_ASCD = X"2F"
						  OR COUNTER_ASCD = X"5D"
						  OR COUNTER_PTX = X"01"
						ELSE '0';
	WR_L			<= '1'
						WHEN COUNTER_ASCD = X"2E"
						ELSE '0';
	RD_PARAMS	<= '1'
						WHEN COUNTER_ASCD = X"33"
						ELSE '0';
	WR_IV			<= '1'
						WHEN (COUNTER_ASCD = X"5C" AND DRL_ASCD = '1')
						  OR COUNTER_ASCD = X"8A"
						ELSE '0';
	DBL_L1		<= '1'
						WHEN COUNTER_ASCD = X"5C"
						ELSE '0';
	RD_ASCD		<= '1'
						WHEN COUNTER_ASCD = X"5F" AND DRL_ASCD = '1'
						ELSE '0';
	RD_PTX		<= '1'
						WHEN DRL_PTX = '1' AND DRL_ASCD = '0' AND COUNTER_PTX = X"03"
						ELSE '0';
	LOAD_IV		<= '1'
						WHEN COUNTER_ASCD = X"5D" OR COUNTER_ASCD = X"8B"
						ELSE '0';
	WR_RO			<= '1'
						WHEN COUNTER_PTX = X"2F"
						ELSE '0';
	DBL_L			<= '1'
						WHEN COUNTER_PTX = X"01"
						ELSE '0';
						
						
	RD_L1			<= '1'
						WHEN COUNTER_ASCD = X"33" OR COUNTER_ASCD = X"61"
						ELSE '0';
	RD_L			<= '1'
						WHEN COUNTER_ASCD = X"FF" --DRL_PTX = '1' AND DRL_ASCD = '0' AND 
						ELSE '0';
	WR_PTX		<= '1'
						WHEN WR = '1' AND ADDR_WR = X"11111111"
						ELSE '0';
	WR_ASCD		<= '1'
						WHEN WR = '1' AND ADDR_WR = X"22222222"
						ELSE '0';
	RD_CTX		<= '1'
						WHEN RD = '1' AND ADDR_WR = X"33333333"
						ELSE '0';
END ARCHITECTURE;