LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY PARAMS_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		RD			:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DATA_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		TAG_INTVL:OUT STD_LOGIC_VECTOR(15 downto 0);
		TAG_LEN	:OUT STD_LOGIC_VECTOR(7 downto 0);
		NPUB		:OUT STD_LOGIC_VECTOR(63 downto 0);
		CONCAT	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE PARAMS_REG_ARCH OF PARAMS_REG IS
	SIGNAL PARAMETERS	:STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			PARAMETERS	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				IF ADDR_WR = X"4" THEN
					PARAMETERS(127 downto 96) <= DATA_WR;
				END IF;
				IF ADDR_WR = X"5" THEN
					PARAMETERS(95 downto 64) <= DATA_WR;
				END IF;
				IF ADDR_WR = X"6" THEN
					PARAMETERS(63 downto 32) <= DATA_WR;
				END IF;
				IF ADDR_WR = X"7" THEN
					PARAMETERS(31 downto 0) <= DATA_WR;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	
	NPUB			<= PARAMETERS(127 downto 64);
	TAG_INTVL	<= PARAMETERS(63 downto 48);
	TAG_LEN		<= PARAMETERS(47 downto 40);
	CONCAT		<= PARAMETERS
						WHEN RD = '1'
						ELSE (OTHERS => '0');
END ARCHITECTURE;