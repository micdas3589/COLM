-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.0 Build 145 04/22/2015 Patches 0.01we SJ Web Edition"
-- CREATED		"Tue Dec 26 22:06:14 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY COLM IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		INIT :  IN  STD_LOGIC;
		WR :  IN  STD_LOGIC;
		RD :  IN  STD_LOGIC;
		ADDR_WR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DIN :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DOUT :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COLM;

ARCHITECTURE bdf_type OF COLM IS 

COMPONENT mem_out
	PORT(CLK : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ascd_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT xor128
	PORT(DIN1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT control
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 DRL_ASCD : IN STD_LOGIC;
		 DRL_PTX : IN STD_LOGIC;
		 DRL_CTX : IN STD_LOGIC;
		 DRL_TAG : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 TAG_CTR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TAG_INTVL : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TAG_LEN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 WR_PTX : OUT STD_LOGIC;
		 WR_ASCD : OUT STD_LOGIC;
		 WR_CTX : OUT STD_LOGIC;
		 WR_TAG : OUT STD_LOGIC;
		 RD_PTX : OUT STD_LOGIC;
		 RD_ASCD : OUT STD_LOGIC;
		 RD_PARAMS : OUT STD_LOGIC;
		 RD_CTX : OUT STD_LOGIC;
		 RD_TAG : OUT STD_LOGIC;
		 WR_L : OUT STD_LOGIC;
		 DBL_L : OUT STD_LOGIC;
		 DBL_L1 : OUT STD_LOGIC;
		 DBL_L2 : OUT STD_LOGIC;
		 WR_IV : OUT STD_LOGIC;
		 RD_L : OUT STD_LOGIC;
		 RD_L1 : OUT STD_LOGIC;
		 WR_RO : OUT STD_LOGIC;
		 LOAD_IV : OUT STD_LOGIC;
		 INIT_EK1 : OUT STD_LOGIC;
		 INIT_EK3 : OUT STD_LOGIC;
		 RUN_EK1 : OUT STD_LOGIC;
		 RUN_EK3 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT mem_out_32
	PORT(CLK : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ctx_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ek
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 RUN : IN STD_LOGIC;
		 KEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_OUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT iv_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 DATA_WR : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 IV : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT key_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 KEY : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT l_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 DBL_L : IN STD_LOGIC;
		 DBL_L1 : IN STD_LOGIC;
		 DBL_L2 : IN STD_LOGIC;
		 RD_L : IN STD_LOGIC;
		 RD_L1 : IN STD_LOGIC;
		 DATA_WR : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 PTX_CTR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 LA : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LB1 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LC2 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or128
	PORT(DIN1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or32
	PORT(DIN1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT params_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 CONCAT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 TAG_INTVL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TAG_LEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ptx_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 PTX_CTR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 TAG_CTR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ro
	PORT(INPUT1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 INPUT2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 OUTPUT1 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 OUTPUT2 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ro_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 LOAD_IV : IN STD_LOGIC;
		 WR_RO : IN STD_LOGIC;
		 IV_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 RO_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 RO : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT tag_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	DBL_L :  STD_LOGIC;
SIGNAL	DBL_L1 :  STD_LOGIC;
SIGNAL	DBL_L2 :  STD_LOGIC;
SIGNAL	DRL_ASCD :  STD_LOGIC;
SIGNAL	DRL_CTX :  STD_LOGIC;
SIGNAL	DRL_PTX :  STD_LOGIC;
SIGNAL	DRL_TAG :  STD_LOGIC;
SIGNAL	INIT_EK1 :  STD_LOGIC;
SIGNAL	INIT_EK3 :  STD_LOGIC;
SIGNAL	IV :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	KEY :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LB1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LC2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LOAD_IV :  STD_LOGIC;
SIGNAL	PTX_CTR :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	RD_ASCD :  STD_LOGIC;
SIGNAL	RD_CTX :  STD_LOGIC;
SIGNAL	RD_L :  STD_LOGIC;
SIGNAL	RD_L1 :  STD_LOGIC;
SIGNAL	RD_PARAMS :  STD_LOGIC;
SIGNAL	RD_PTX :  STD_LOGIC;
SIGNAL	RD_TAG :  STD_LOGIC;
SIGNAL	RO_IN :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	RO_OUT :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	RUN_EK1 :  STD_LOGIC;
SIGNAL	RUN_EK3 :  STD_LOGIC;
SIGNAL	STATE_IN1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_IN3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUTA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUTB :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUTC :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	TAG_CTR :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	TAG_INTVL :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	TAG_LEN :  STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL	WR_ASCD :  STD_LOGIC;
SIGNAL	WR_CTX :  STD_LOGIC;
SIGNAL	WR_IV :  STD_LOGIC;
SIGNAL	WR_L :  STD_LOGIC;
SIGNAL	WR_PTX :  STD_LOGIC;
SIGNAL	WR_RO :  STD_LOGIC;
SIGNAL	WR_TAG :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC_VECTOR(127 DOWNTO 0);


BEGIN 



b2v_ASCD_MEM_OUT : mem_out
PORT MAP(CLK => CLK,
		 LOAD => RD_ASCD,
		 DIN => SYNTHESIZED_WIRE_0,
		 DOUT => SYNTHESIZED_WIRE_9);


b2v_ASCD_MEMORY : ascd_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_ASCD,
		 LOAD => RD_ASCD,
		 DIN => DIN,
		 DRL => DRL_ASCD,
		 DOUT => SYNTHESIZED_WIRE_0);


b2v_ASCD_XOR : xor128
PORT MAP(DIN1 => LB1,
		 DIN2 => SYNTHESIZED_WIRE_1,
		 DOUT => SYNTHESIZED_WIRE_5);


b2v_CONTROL : control
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 RD => RD,
		 DRL_ASCD => DRL_ASCD,
		 DRL_PTX => DRL_PTX,
		 DRL_CTX => DRL_CTX,
		 DRL_TAG => DRL_TAG,
		 ADDR_WR => ADDR_WR,
		 TAG_CTR => TAG_CTR,
		 TAG_INTVL => TAG_INTVL,
		 TAG_LEN => TAG_LEN,
		 WR_PTX => WR_PTX,
		 WR_ASCD => WR_ASCD,
		 WR_CTX => WR_CTX,
		 WR_TAG => WR_TAG,
		 RD_PTX => RD_PTX,
		 RD_ASCD => RD_ASCD,
		 RD_PARAMS => RD_PARAMS,
		 RD_CTX => RD_CTX,
		 RD_TAG => RD_TAG,
		 WR_L => WR_L,
		 DBL_L => DBL_L,
		 DBL_L1 => DBL_L1,
		 DBL_L2 => DBL_L2,
		 WR_IV => WR_IV,
		 RD_L => RD_L,
		 RD_L1 => RD_L1,
		 WR_RO => WR_RO,
		 LOAD_IV => LOAD_IV,
		 INIT_EK1 => INIT_EK1,
		 INIT_EK3 => INIT_EK3,
		 RUN_EK1 => RUN_EK1,
		 RUN_EK3 => RUN_EK3);


b2v_CTX_MEM_OUT : mem_out_32
PORT MAP(CLK => CLK,
		 LOAD => RD_CTX,
		 DIN => SYNTHESIZED_WIRE_2,
		 DOUT => SYNTHESIZED_WIRE_6);


b2v_CTX_MEMORY : ctx_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_CTX,
		 LOAD => RD_CTX,
		 DIN => SYNTHESIZED_WIRE_3,
		 DRL => DRL_CTX,
		 DOUT => SYNTHESIZED_WIRE_2);


b2v_EK1 : ek
PORT MAP(CLK => CLK,
		 INIT => INIT_EK1,
		 RUN => RUN_EK1,
		 KEY => KEY,
		 STATE_IN => STATE_IN1,
		 STATE_OUT => STATE_OUTA);


b2v_EK2 : ek
PORT MAP(CLK => CLK,
		 INIT => INIT_EK3,
		 RUN => RUN_EK3,
		 KEY => KEY,
		 STATE_IN => RO_IN,
		 STATE_OUT => STATE_OUTB);


b2v_EK2_XOR3 : xor128
PORT MAP(DIN1 => STATE_OUTB,
		 DIN2 => LC2,
		 DOUT => SYNTHESIZED_WIRE_13);


b2v_EK3 : ek
PORT MAP(CLK => CLK,
		 INIT => INIT_EK3,
		 RUN => RUN_EK3,
		 KEY => KEY,
		 STATE_IN => STATE_IN3,
		 STATE_OUT => STATE_OUTC);


b2v_EK3_XOR : xor128
PORT MAP(DIN1 => STATE_OUTC,
		 DIN2 => LC2,
		 DOUT => SYNTHESIZED_WIRE_3);


b2v_IV_REG : iv_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR_IV,
		 DATA_WR => STATE_OUTA,
		 IV => IV);


b2v_KEY_REG : key_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 KEY => KEY);


b2v_L_REG : l_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR_L,
		 DBL_L => DBL_L,
		 DBL_L1 => DBL_L1,
		 DBL_L2 => DBL_L2,
		 RD_L => RD_L,
		 RD_L1 => RD_L1,
		 DATA_WR => STATE_OUTA,
		 PTX_CTR => PTX_CTR,
		 LA => LA,
		 LB1 => LB1,
		 LC2 => LC2);


b2v_OR : or128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_4,
		 DIN2 => SYNTHESIZED_WIRE_5,
		 DOUT => STATE_IN1);


b2v_OR32 : or32
PORT MAP(DIN1 => SYNTHESIZED_WIRE_6,
		 DIN2 => SYNTHESIZED_WIRE_7,
		 DOUT => DOUT);


b2v_PARAMS_OR : or128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_8,
		 DIN2 => SYNTHESIZED_WIRE_9,
		 DOUT => SYNTHESIZED_WIRE_1);


b2v_PARAMS_REG : params_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 RD => RD_PARAMS,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 CONCAT => SYNTHESIZED_WIRE_8,
		 TAG_INTVL => TAG_INTVL,
		 TAG_LEN => TAG_LEN);


b2v_PTX_MEM_OUT : mem_out
PORT MAP(CLK => CLK,
		 LOAD => RD_PTX,
		 DIN => SYNTHESIZED_WIRE_10,
		 DOUT => SYNTHESIZED_WIRE_11);


b2v_PTX_MEMORY : ptx_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_PTX,
		 LOAD => RD_PTX,
		 DIN => DIN,
		 DRL => DRL_PTX,
		 DOUT => SYNTHESIZED_WIRE_10,
		 PTX_CTR => PTX_CTR,
		 TAG_CTR => TAG_CTR);


b2v_PTX_XOR : xor128
PORT MAP(DIN1 => LA,
		 DIN2 => SYNTHESIZED_WIRE_11,
		 DOUT => SYNTHESIZED_WIRE_4);


b2v_RO : ro
PORT MAP(INPUT1 => STATE_OUTA,
		 INPUT2 => RO_OUT,
		 OUTPUT1 => STATE_IN3,
		 OUTPUT2 => RO_IN);


b2v_RO_REG : ro_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 LOAD_IV => LOAD_IV,
		 WR_RO => WR_RO,
		 IV_IN => IV,
		 RO_IN => RO_IN,
		 RO => RO_OUT);


b2v_TAG_MEM_OUT : mem_out_32
PORT MAP(CLK => CLK,
		 LOAD => RD_TAG,
		 DIN => SYNTHESIZED_WIRE_12,
		 DOUT => SYNTHESIZED_WIRE_7);


b2v_TAG_MEMORY : tag_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_TAG,
		 LOAD => RD_TAG,
		 DIN => SYNTHESIZED_WIRE_13,
		 DRL => DRL_TAG,
		 DOUT => SYNTHESIZED_WIRE_12);


END bdf_type;