LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY RO IS
	PORT (
		INPUT1	:IN STD_LOGIC_VECTOR(127 downto 0);
		INPUT2	:IN STD_LOGIC_VECTOR(127 downto 0);
		OUTPUT1	:OUT STD_LOGIC_VECTOR(127 downto 0);
		OUTPUT2	:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE RO_ARCH OF RO IS
BEGIN
	OUTPUT1	<= INPUT1 XOR INPUT2 XOR ('0' & INPUT2(126 downto 0)) XOR X"87" --multiply by 3
					WHEN INPUT2(127) = '1' ELSE
					INPUT1 XOR INPUT2 XOR ('0' & INPUT2(126 downto 0));
	OUTPUT2	<= INPUT1 XOR ('0' & INPUT2(126 downto 0)) XOR X"87" -- multiply by 2
					WHEN INPUT2(127) = '1' ELSE
					INPUT1 XOR ('0' & INPUT2(126 downto 0));
END ARCHITECTURE;