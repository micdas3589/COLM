 LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY PTX_TAG_GENERATOR IS
	PORT (
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		ADDR_WR	:IN STD_LOGIC_VECTOR(31 downto 0);
		DIN		:IN STD_LOGIC_VECTOR(31 downto 0);

		PTX_TAG	:OUT STD_LOGIC_VECTOR(31 downto 0)
	);
END ENTITY;

ARCHITECTURE ARCH_PTX_TAG_GENERATOR OF PTX_TAG_GENERATOR IS
	SIGNAL PTX_CTR			:STD_LOGIC_VECTOR(1 downto 0);
	SIGNAL PTX_TAG_VAL	:STD_LOGIC_VECTOR(127 downto 0);
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			PTX_CTR		<= (OTHERS => '0');
			PTX_TAG_VAL	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' AND ADDR_WR = X"11111111" THEN
				IF PTX_CTR = "00" THEN
					PTX_TAG_VAL(127 downto 96)	<= PTX_TAG_VAL(127 downto 96) XOR DIN;
				END IF;
				IF PTX_CTR = "01" THEN
					PTX_TAG_VAL(95 downto 64)	<= PTX_TAG_VAL(95 downto 64) XOR DIN;
				END IF;
				IF PTX_CTR = "10" THEN
					PTX_TAG_VAL(63 downto 32)	<= PTX_TAG_VAL(63 downto 32) XOR DIN;
				END IF;
				IF PTX_CTR = "11" THEN
					PTX_TAG_VAL(31 downto 0)	<= PTX_TAG_VAL(31 downto 0) XOR DIN;
				END IF;
				
				PTX_CTR	<= PTX_CTR + 1;
			END IF;
			
			IF WR = '1' AND ADDR_WR = X"55555555" THEN
				PTX_CTR	<= PTX_CTR + 1;
			END IF;
		END IF;
	END PROCESS;
	
	PTX_TAG	<=  PTX_TAG_VAL(127 downto 96)
			  WHEN PTX_CTR = "00" AND WR = '1' AND ADDR_WR = X"55555555"
			  ELSE PTX_TAG_VAL(95 downto 64)
			  WHEN PTX_CTR = "01" AND WR = '1' AND ADDR_WR = X"55555555"
			  ELSE PTX_TAG_VAL(63 downto 32)
			  WHEN PTX_CTR = "10" AND WR = '1' AND ADDR_WR = X"55555555"
			  ELSE PTX_TAG_VAL(31 downto 0)
			  WHEN PTX_CTR = "11" AND WR = '1' AND ADDR_WR = X"55555555"
			  ELSE (OTHERS => '0');
END ARCHITECTURE;