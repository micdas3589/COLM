LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY IV_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		RD			:IN STD_LOGIC;
		DATA_WR	:IN STD_LOGIC_VECTOR(127 downto 0);
		IV			:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE IV_REG_ARCH OF IV_REG IS
	SIGNAL STATE	:STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			STATE	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				STATE	<= STATE XOR DATA_WR;
			END IF;
		END IF;
	END PROCESS;
	
	IV	<= STATE
			WHEN RD = '1'
			ELSE (OTHERS => '0');
END ARCHITECTURE;