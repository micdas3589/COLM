LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RO_REG IS
	PORT
	(
		CLK	:IN STD_LOGIC;
		INIT	:IN STD_LOGIC;
		WR		:IN STD_LOGIC;
		RO_IN	:IN STD_LOGIC_VECTOR(127 downto 0);
		RO		:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE RO_REG_ARCH OF RO_REG IS
	SIGNAL RO_STATE	:STD_LOGIC_VECTOR(127 downto 0);
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			RO_STATE	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				RO_STATE	<= RO_IN;
			END IF;
		END IF;
		
		RO	<= RO_STATE;
	END PROCESS;
END ARCHITECTURE;