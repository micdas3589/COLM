LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.NUMERIC_STD.ALL;

ENTITY L_REG_TB IS END ENTITY;

ARCHITECTURE ARCH_L_REG_TB OF L_REG_TB IS
	COMPONENT L_REG IS PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		DATA_WR	:IN STD_LOGIC_VECTOR(127 downto 0);
		DBL_L		:IN STD_LOGIC;
		DBL_L1	:IN STD_LOGIC;
		DBL_L2	:IN STD_LOGIC;
		RD_L		:IN STD_LOGIC;
		RD_L1		:IN STD_LOGIC;
		PTX_CTR	:IN STD_LOGIC_VECTOR(7 downto 0);
		LA			:OUT STD_LOGIC_VECTOR(127 downto 0);
		LB1		:OUT STD_LOGIC_VECTOR(127 downto 0);
		LC2		:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
	END COMPONENT;

	SIGNAL CLK		: STD_LOGIC := '0';
	SIGNAL INIT		: STD_LOGIC := '0';
	SIGNAL WR			: STD_LOGIC := '0';
	SIGNAL DATA_WR	: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL DBL_L		: STD_LOGIC := '0';
	SIGNAL DBL_L1	: STD_LOGIC := '0';
	SIGNAL DBL_L2	: STD_LOGIC := '0';
	SIGNAL RD_L		: STD_LOGIC := '0';
	SIGNAL RD_L1		: STD_LOGIC := '0';
	SIGNAL PTX_CTR	: STD_LOGIC_VECTOR(7 downto 0);
	SIGNAL LA			: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL LB1		: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL LC2		: STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	
	SIGNAL CLKp :time := 40 ns;
BEGIN
	tb: L_REG PORT MAP (CLK, INIT, WR, DATA_WR, DBL_L, DBL_L1, DBL_L2, RD_L, RD_L1, PTX_CTR, LA, LB1, LC2);

	PROCESS
	BEGIN
		CLK <= '0'; wait for CLKp / 2;
		CLK <= '1'; wait for CLKp / 2;
	END PROCESS;

	PROCESS
	BEGIN
		INIT <= '1'; WR <= '0'; DATA_WR <= X"00000000000000000000000000000000"; DBL_L <= '1'; DBL_L1 <= '1'; DBL_L2 <= '1'; RD_L <= '1'; RD_L1 <= '1'; PTX_CTR <= X"00"; wait for CLKp;
		INIT <= '0'; WR <= '1'; DATA_WR <= X"11111111111111111111111111111111"; DBL_L <= '1'; DBL_L1 <= '1'; DBL_L2 <= '1'; RD_L <= '1'; RD_L1 <= '1'; PTX_CTR <= X"00"; wait for CLKp;
		INIT <= '0'; WR <= '0'; DATA_WR <= X"22222222222222222222222222222222"; DBL_L <= '1'; DBL_L1 <= '1'; DBL_L2 <= '1'; RD_L <= '1'; RD_L1 <= '1'; PTX_CTR <= X"00"; wait for CLKp;
		INIT <= '0'; WR <= '1'; DATA_WR <= X"00000000000000000000000000000000"; DBL_L <= '1'; DBL_L1 <= '1'; DBL_L2 <= '1'; RD_L <= '1'; RD_L1 <= '1'; PTX_CTR <= X"00"; wait for 10*CLKp;
		wait;
	END PROCESS;
END ARCHITECTURE;