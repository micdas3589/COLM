LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MAX_ADDR_REG IS
	PORT
	(
		CLK			:IN STD_LOGIC;
		INIT			:IN STD_LOGIC;
		INCR_PTX		:IN STD_LOGIC;
		INCR_ASCD	:IN STD_LOGIC;
		MAX_PTX		:OUT STD_LOGIC_VECTOR(7 downto 0);
		MAX_ASCD		:OUT STD_LOGIC_VECTOR(7 downto 0)
	);
END ENTITY;

ARCHITECTURE MAX_ADDR_REG_ARCH OF MAX_ADDR_REG IS
	SIGNAL PTX_MAX_ADDR	:STD_LOGIC_VECTOR(7 downto 0) := (OTHERS => '0');
	SIGNAL ASCD_MAX_ADDR	:STD_LOGIC_VECTOR(7 downto 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			PTX_MAX_ADDR	<= X"0";
			ASCD_MAX_ADDR	<= X"100";
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF INCR_PTX = '1' THEN
				PTX_MAX_ADDR	<= PTX_MAX_ADDR + 1;
			END IF;
			IF INCR_ASCD = '1' THEN
				ASCD_MAX_ADDR	<= ASCD_MAX_ADDR + 1;
			END IF;
		END IF;
	END PROCESS;
	
	MAX_PTX	<= PTX_MAX_ADDR;
	MAX_ASCD	<= ASCD_MAX_ADDR;
END ARCHITECTURE;