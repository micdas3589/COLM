-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.0 Build 145 04/22/2015 Patches 0.01we SJ Web Edition"
-- CREATED		"Tue Aug 08 20:22:35 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY COLM IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		INIT :  IN  STD_LOGIC;
		WR :  IN  STD_LOGIC;
		ADDR_WR :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DIN :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		DOUT :  OUT  STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COLM;

ARCHITECTURE bdf_type OF COLM IS 

COMPONENT control
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 DRL_ASCD : IN STD_LOGIC;
		 DRL_PTX : IN STD_LOGIC;
		 DRL_CTX : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 WR_PTX : OUT STD_LOGIC;
		 WR_ASCD : OUT STD_LOGIC;
		 WR_CTX : OUT STD_LOGIC;
		 RD_PTX : OUT STD_LOGIC;
		 RD_ASCD : OUT STD_LOGIC;
		 RD_PARAMS : OUT STD_LOGIC;
		 RD_CTX : OUT STD_LOGIC;
		 WR_L : OUT STD_LOGIC;
		 DBL_L : OUT STD_LOGIC;
		 DBL_L1 : OUT STD_LOGIC;
		 DBL_L2 : OUT STD_LOGIC;
		 WR_IV : OUT STD_LOGIC;
		 RD_IV : OUT STD_LOGIC;
		 RD_L : OUT STD_LOGIC;
		 RD_L1 : OUT STD_LOGIC;
		 WR_RO : OUT STD_LOGIC;
		 INIT_EK1 : OUT STD_LOGIC;
		 INIT_EK2 : OUT STD_LOGIC;
		 INIT_EK3 : OUT STD_LOGIC;
		 RUN_EK1 : OUT STD_LOGIC;
		 RUN_EK2 : OUT STD_LOGIC;
		 RUN_EK3 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT l_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 DBL_L : IN STD_LOGIC;
		 DBL_L1 : IN STD_LOGIC;
		 DBL_L2 : IN STD_LOGIC;
		 RD_L : IN STD_LOGIC;
		 RD_L1 : IN STD_LOGIC;
		 DATA_WR : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LA : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LB1 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 LC2 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ek
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 RUN : IN STD_LOGIC;
		 KEY : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_IN : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 STATE_OUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT iv_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 DATA_WR : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 IV : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT key_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 KEY : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT params_reg
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 WR : IN STD_LOGIC;
		 RD : IN STD_LOGIC;
		 ADDR_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_WR : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 CONCAT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
		 NPUB : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
		 TAG_INTVL : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 TAG_LEN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ascd_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ptx_memory
	PORT(CLK : IN STD_LOGIC;
		 INIT : IN STD_LOGIC;
		 STORE : IN STD_LOGIC;
		 LOAD : IN STD_LOGIC;
		 DIN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DRL : OUT STD_LOGIC;
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT xor128
	PORT(DIN1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

COMPONENT or128
	PORT(DIN1 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DIN2 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		 DOUT : OUT STD_LOGIC_VECTOR(127 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	DATA_WR :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	DBL_L :  STD_LOGIC;
SIGNAL	DBL_L1 :  STD_LOGIC;
SIGNAL	DBL_L2 :  STD_LOGIC;
SIGNAL	DRL_ASCD :  STD_LOGIC;
SIGNAL	DRL_CTX :  STD_LOGIC;
SIGNAL	DRL_PTX :  STD_LOGIC;
SIGNAL	INIT_EK1 :  STD_LOGIC;
SIGNAL	IV :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	KEY :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LA :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LB1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	LC2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	RD :  STD_LOGIC;
SIGNAL	RD_ASCD :  STD_LOGIC;
SIGNAL	RD_IV :  STD_LOGIC;
SIGNAL	RD_L :  STD_LOGIC;
SIGNAL	RD_L1 :  STD_LOGIC;
SIGNAL	RD_PARAMS :  STD_LOGIC;
SIGNAL	RD_PTX :  STD_LOGIC;
SIGNAL	RUN_EK1 :  STD_LOGIC;
SIGNAL	STATE_IN :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	STATE_OUT :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	WR_ASCD :  STD_LOGIC;
SIGNAL	WR_IV :  STD_LOGIC;
SIGNAL	WR_PTX :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(127 DOWNTO 0);


BEGIN 



b2v_inst : control
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 RD => RD,
		 DRL_ASCD => DRL_ASCD,
		 DRL_PTX => DRL_PTX,
		 DRL_CTX => DRL_CTX,
		 ADDR_WR => ADDR_WR,
		 WR_PTX => WR_PTX,
		 WR_ASCD => WR_ASCD,
		 RD_PTX => RD_PTX,
		 RD_ASCD => RD_ASCD,
		 RD_PARAMS => RD_PARAMS,
		 DBL_L => DBL_L,
		 DBL_L1 => DBL_L1,
		 DBL_L2 => DBL_L2,
		 RD_IV => RD_IV,
		 RD_L => RD_L,
		 RD_L1 => RD_L1,
		 INIT_EK1 => INIT_EK1,
		 RUN_EK1 => RUN_EK1);


b2v_inst10 : l_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 DBL_L => DBL_L,
		 DBL_L1 => DBL_L1,
		 DBL_L2 => DBL_L2,
		 RD_L => RD_L,
		 RD_L1 => RD_L1,
		 DATA_WR => DATA_WR,
		 LA => LA,
		 LB1 => LB1);


b2v_inst11 : ek
PORT MAP(CLK => CLK,
		 INIT => INIT_EK1,
		 RUN => RUN_EK1,
		 KEY => KEY,
		 STATE_IN => STATE_IN,
		 STATE_OUT => STATE_OUT);


b2v_inst13 : iv_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR_IV,
		 RD => RD_IV,
		 DATA_WR => STATE_OUT);


b2v_inst14 : key_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 KEY => KEY);


b2v_inst2 : params_reg
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 WR => WR,
		 RD => RD_PARAMS,
		 ADDR_WR => ADDR_WR,
		 DATA_WR => DIN,
		 CONCAT => SYNTHESIZED_WIRE_2);


b2v_inst3 : ascd_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_ASCD,
		 LOAD => RD_ASCD,
		 DIN => DIN,
		 DRL => DRL_ASCD,
		 DOUT => SYNTHESIZED_WIRE_3);


b2v_inst4 : ptx_memory
PORT MAP(CLK => CLK,
		 INIT => INIT,
		 STORE => WR_PTX,
		 LOAD => RD_PTX,
		 DIN => DIN,
		 DRL => DRL_PTX,
		 DOUT => SYNTHESIZED_WIRE_1);


b2v_inst5 : xor128
PORT MAP(DIN1 => LB1,
		 DIN2 => SYNTHESIZED_WIRE_0,
		 DOUT => SYNTHESIZED_WIRE_5);


b2v_inst6 : xor128
PORT MAP(DIN1 => LA,
		 DIN2 => SYNTHESIZED_WIRE_1,
		 DOUT => SYNTHESIZED_WIRE_4);


b2v_inst8 : or128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_2,
		 DIN2 => SYNTHESIZED_WIRE_3,
		 DOUT => SYNTHESIZED_WIRE_0);


b2v_inst9 : or128
PORT MAP(DIN1 => SYNTHESIZED_WIRE_4,
		 DIN2 => SYNTHESIZED_WIRE_5,
		 DOUT => STATE_IN);

DOUT <= STATE_OUT;

END bdf_type;