LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY L_REG IS
	PORT
	(
		CLK		:IN STD_LOGIC;
		INIT		:IN STD_LOGIC;
		WR			:IN STD_LOGIC;
		DATA_WR	:IN STD_LOGIC_VECTOR(127 downto 0);
		L			:OUT STD_LOGIC_VECTOR(127 downto 0);
		L1			:OUT STD_LOGIC_VECTOR(127 downto 0);
		L2			:OUT STD_LOGIC_VECTOR(127 downto 0)
	);
END ENTITY;

ARCHITECTURE L_REG_ARCH OF L_REG IS
	SIGNAL COUNTER	:STD_LOGIC_VECTOR(2 downto 0) := (OTHERS => '0');
	SIGNAL L_VALUE	:STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
	SIGNAL L2_VALUE	:STD_LOGIC_VECTOR(127 downto 0) := (OTHERS => '0');
BEGIN
	PROCESS(CLK, INIT)
	BEGIN
		IF INIT = '1' THEN
			COUNTER	<= (OTHERS => '0');
			L_VALUE	<= (OTHERS => '0');
		ELSIF CLK = '1' AND CLK'EVENT THEN
			IF WR = '1' THEN
				L_VALUE	<= DATA_WR;
				L2_VALUE	<= DATA_WR;
				COUNTER	<= COUNTER + 1;
			END IF;
			IF COUNTER = X"1" OR COUNTER = X"2" THEN
				IF L2_VALUE(127) = '1' THEN
					L2_VALUE	<= L2_VALUE XOR ('0' & L2_VALUE(126 downto 0)) XOR X"87";
				ELSE
					L2_VALUE	<= L2_VALUE XOR ('0' & L2_VALUE(126 downto 0));
				END IF;
				
				COUNTER	<= COUNTER + 1;
			END IF;
		END IF;
	END PROCESS;
	
	L	<= L_VALUE;
	L1	<= L_VALUE XOR ('0' & L_VALUE(126 downto 0)) XOR X"87"
			WHEN L_VALUE(127) = '1' ELSE
			L_VALUE XOR ('0' & L_VALUE(126 downto 0));
	L2	<= L2_VALUE;
END ARCHITECTURE;